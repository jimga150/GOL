----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:12:33 01/21/2019 
-- Design Name: 
-- Module Name:    SegmentReaderSM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SegmentReaderSM is
    Port ( start_read, rd_empty : in  STD_LOGIC;
           col_plus_one : in  STD_LOGIC_VECTOR (7 downto 0);
           segment : in  STD_LOGIC_VECTOR (7 downto 0);
           done, rd_en, img_src_en : out  STD_LOGIC;
           col : out  STD_LOGIC_VECTOR (7 downto 0));
end SegmentReaderSM;

architecture Behavioral of SegmentReaderSM is

begin


end Behavioral;

